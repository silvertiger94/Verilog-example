`timescale 1ns / 1ns
`include "macro.svh"
